`timescale 1ns/1ps
//////////////////////////////////////////////////////////////////////////////////
//  
//  
// Code by : Sananda Ghosh, Amogh Halgeri from Upenn
//
// Date:   06/29/2011 - modified July 13 2012 (Madhura)
// Module Name:    trial128bit.v
//  
// Description: The 128 bit strip data is analyzed and more than two hits occur, they are ignored.
//		The location of the hits are denoted by a 7 bit address, and the one adjacent bit is used to denote the
//		presence of a second consecutive hit.
//
//////////////////////////////////////////////////////////////////////////////////

module trial128bit(single,double,totaladdr);
reg [127:0]data;
input [127:0]single;
input [127:0]double;
//input BCclk;
output [15:0]totaladdr;			
//output count;
wire [7:0] first,second,third;

//reg count;
wire [6:0] firsttemp;
wire [127:0] mask;
reg [127:0] datatemp;
wire lclClk;


   always@(single or double or mask)
     begin
	datatemp <= mask & (single | double);
	
     end
   
   
   
   //This gives the first hit cluster location 
   assign first = 	(single[0])? {1'b0,7'd0} : (double[0]) ? {1'b1,7'd0} :
		  (single[1])? {1'b0,7'd1} : (double[1]) ? {1'b1,7'd1} :
		  (single[2])? {1'b0,7'd2} : (double[2]) ? {1'b1,7'd2} :
		  (single[3])? {1'b0,7'd3} : (double[3]) ? {1'b1,7'd3} :
		  (single[4])? {1'b0,7'd4} : (double[4]) ? {1'b1,7'd4} :
		  (single[5])? {1'b0,7'd5} : (double[5]) ? {1'b1,7'd5} :
		  (single[6])? {1'b0,7'd6} : (double[6]) ? {1'b1,7'd6} :
		  (single[7])? {1'b0,7'd7} : (double[7]) ? {1'b1,7'd7} :
		  (single[8])? {1'b0,7'd8} : (double[8]) ? {1'b1,7'd8} :
		  (single[9])? {1'b0,7'd9} : (double[9]) ? {1'b1,7'd9} :
		  (single[10])? {1'b0,7'd10} : (double[10]) ? {1'b1,7'd10} :
		  (single[11])? {1'b0,7'd11} : (double[11]) ? {1'b1,7'd11} :
		  (single[12])? {1'b0,7'd12} : (double[12]) ? {1'b1,7'd12} :
		  (single[13])? {1'b0,7'd13} : (double[13]) ? {1'b1,7'd13} :
		  (single[14])? {1'b0,7'd14} : (double[14]) ? {1'b1,7'd14} :
		  (single[15])? {1'b0,7'd15} : (double[15]) ? {1'b1,7'd15} :
		  (single[16])? {1'b0,7'd16} : (double[16]) ? {1'b1,7'd16} :
		  (single[17])? {1'b0,7'd17} : (double[17]) ? {1'b1,7'd17} :
		  (single[18])? {1'b0,7'd18} : (double[18]) ? {1'b1,7'd18} :
		  (single[19])? {1'b0,7'd19} : (double[19]) ? {1'b1,7'd19} :
		  (single[20])? {1'b0,7'd20} : (double[20]) ? {1'b1,7'd20} :
		  (single[21])? {1'b0,7'd21} : (double[21]) ? {1'b1,7'd21} :
		  (single[22])? {1'b0,7'd22} : (double[22]) ? {1'b1,7'd22} :
		  (single[23])? {1'b0,7'd23} : (double[23]) ? {1'b1,7'd23} :
		  (single[24])? {1'b0,7'd24} : (double[24]) ? {1'b1,7'd24} :
		  (single[25])? {1'b0,7'd25} : (double[25]) ? {1'b1,7'd25} :
		  (single[26])? {1'b0,7'd26} : (double[26]) ? {1'b1,7'd26} :
		  (single[27])? {1'b0,7'd27} : (double[27]) ? {1'b1,7'd27} :
		  (single[28])? {1'b0,7'd28} : (double[28]) ? {1'b1,7'd28} :
		  (single[29])? {1'b0,7'd29} : (double[29]) ? {1'b1,7'd29} :
		  (single[30])? {1'b0,7'd30} : (double[30]) ? {1'b1,7'd30} :
		  (single[31])? {1'b0,7'd31} : (double[31]) ? {1'b1,7'd31} :
		  (single[32])? {1'b0,7'd32} : (double[32]) ? {1'b1,7'd32} :
		  (single[33])? {1'b0,7'd33} : (double[33]) ? {1'b1,7'd33} :
		  (single[34])? {1'b0,7'd34} : (double[34]) ? {1'b1,7'd34} :
		  (single[35])? {1'b0,7'd35} : (double[35]) ? {1'b1,7'd35} :
		  (single[36])? {1'b0,7'd36} : (double[36]) ? {1'b1,7'd36} :
		  (single[37])? {1'b0,7'd37} : (double[37]) ? {1'b1,7'd37} :
		  (single[38])? {1'b0,7'd38} : (double[38]) ? {1'b1,7'd38} :
		  (single[39])? {1'b0,7'd39} : (double[39]) ? {1'b1,7'd39} :
		  (single[40])? {1'b0,7'd40} : (double[40]) ? {1'b1,7'd40} :
		  (single[41])? {1'b0,7'd41} : (double[41]) ? {1'b1,7'd41} :
		  (single[42])? {1'b0,7'd42} : (double[42]) ? {1'b1,7'd42} :
		  (single[43])? {1'b0,7'd43} : (double[43]) ? {1'b1,7'd43} :
		  (single[44])? {1'b0,7'd44} : (double[44]) ? {1'b1,7'd44} :
		  (single[45])? {1'b0,7'd45} : (double[45]) ? {1'b1,7'd45} :
		  (single[46])? {1'b0,7'd46} : (double[46]) ? {1'b1,7'd46} :
		  (single[47])? {1'b0,7'd47} : (double[47]) ? {1'b1,7'd47} :
		  (single[48])? {1'b0,7'd48} : (double[48]) ? {1'b1,7'd48} :
		  (single[49])? {1'b0,7'd49} : (double[49]) ? {1'b1,7'd49} :
		  (single[50])? {1'b0,7'd50} : (double[50]) ? {1'b1,7'd50} :
		  (single[51])? {1'b0,7'd51} : (double[51]) ? {1'b1,7'd51} :
		  (single[52])? {1'b0,7'd52} : (double[52]) ? {1'b1,7'd52} :
		  (single[53])? {1'b0,7'd53} : (double[53]) ? {1'b1,7'd53} :
		  (single[54])? {1'b0,7'd54} : (double[54]) ? {1'b1,7'd54} :
		  (single[55])? {1'b0,7'd55} : (double[55]) ? {1'b1,7'd55} :
		  (single[56])? {1'b0,7'd56} : (double[56]) ? {1'b1,7'd56} :
		  (single[57])? {1'b0,7'd57} : (double[57]) ? {1'b1,7'd57} :
		  (single[58])? {1'b0,7'd58} : (double[58]) ? {1'b1,7'd58} :
		  (single[59])? {1'b0,7'd59} : (double[59]) ? {1'b1,7'd59} :
		  (single[60])? {1'b0,7'd60} : (double[60]) ? {1'b1,7'd60} :
		  (single[61])? {1'b0,7'd61} : (double[61]) ? {1'b1,7'd61} :
		  (single[62])? {1'b0,7'd62} : (double[62]) ? {1'b1,7'd62} :
		  (single[63])? {1'b0,7'd63} : (double[63]) ? {1'b1,7'd63} :
		  (single[64])? {1'b0,7'd64} : (double[64]) ? {1'b1,7'd64} :
		  (single[65])? {1'b0,7'd65} : (double[65]) ? {1'b1,7'd65} :
		  (single[66])? {1'b0,7'd66} : (double[66]) ? {1'b1,7'd66} :
		  (single[67])? {1'b0,7'd67} : (double[67]) ? {1'b1,7'd67} :
		  (single[68])? {1'b0,7'd68} : (double[68]) ? {1'b1,7'd68} :
		  (single[69])? {1'b0,7'd69} : (double[69]) ? {1'b1,7'd69} :
		  (single[70])? {1'b0,7'd70} : (double[70]) ? {1'b1,7'd70} :
		  (single[71])? {1'b0,7'd71} : (double[71]) ? {1'b1,7'd71} :
		  (single[72])? {1'b0,7'd72} : (double[72]) ? {1'b1,7'd72} :
		  (single[73])? {1'b0,7'd73} : (double[73]) ? {1'b1,7'd73} :
		  (single[74])? {1'b0,7'd74} : (double[74]) ? {1'b1,7'd74} :
		  (single[75])? {1'b0,7'd75} : (double[75]) ? {1'b1,7'd75} :
		  (single[76])? {1'b0,7'd76} : (double[76]) ? {1'b1,7'd76} :
		  (single[77])? {1'b0,7'd77} : (double[77]) ? {1'b1,7'd77} :
		  (single[78])? {1'b0,7'd78} : (double[78]) ? {1'b1,7'd78} :
		  (single[79])? {1'b0,7'd79} : (double[79]) ? {1'b1,7'd79} :
		  (single[80])? {1'b0,7'd80} : (double[80]) ? {1'b1,7'd80} :
		  (single[81])? {1'b0,7'd81} : (double[81]) ? {1'b1,7'd81} :
		  (single[82])? {1'b0,7'd82} : (double[82]) ? {1'b1,7'd82} :
		  (single[83])? {1'b0,7'd83} : (double[83]) ? {1'b1,7'd83} :
		  (single[84])? {1'b0,7'd84} : (double[84]) ? {1'b1,7'd84} :
		  (single[85])? {1'b0,7'd85} : (double[85]) ? {1'b1,7'd85} :
		  (single[86])? {1'b0,7'd86} : (double[86]) ? {1'b1,7'd86} :
		  (single[87])? {1'b0,7'd87} : (double[87]) ? {1'b1,7'd87} :
		  (single[88])? {1'b0,7'd88} : (double[88]) ? {1'b1,7'd88} :
		  (single[89])? {1'b0,7'd89} : (double[89]) ? {1'b1,7'd89} :
		  (single[90])? {1'b0,7'd90} : (double[90]) ? {1'b1,7'd90} :
		  (single[91])? {1'b0,7'd91} : (double[91]) ? {1'b1,7'd91} :
		  (single[92])? {1'b0,7'd92} : (double[92]) ? {1'b1,7'd92} :
		  (single[93])? {1'b0,7'd93} : (double[93]) ? {1'b1,7'd93} :
		  (single[94])? {1'b0,7'd94} : (double[94]) ? {1'b1,7'd94} :
		  (single[95])? {1'b0,7'd95} : (double[95]) ? {1'b1,7'd95} :
		  (single[96])? {1'b0,7'd96} : (double[96]) ? {1'b1,7'd96} :
		  (single[97])? {1'b0,7'd97} : (double[97]) ? {1'b1,7'd97} :
		  (single[98])? {1'b0,7'd98} : (double[98]) ? {1'b1,7'd98} :
		  (single[99])? {1'b0,7'd99} : (double[99]) ? {1'b1,7'd99} :
		  (single[100])? {1'b0,7'd100} : (double[100]) ? {1'b1,7'd100} :
		  (single[101])? {1'b0,7'd101} : (double[101]) ? {1'b1,7'd101} :
		  (single[102])? {1'b0,7'd102} : (double[102]) ? {1'b1,7'd102} :
		  (single[103])? {1'b0,7'd103} : (double[103]) ? {1'b1,7'd103} :
		  (single[104])? {1'b0,7'd104} : (double[104]) ? {1'b1,7'd104} :
		  (single[105])? {1'b0,7'd105} : (double[105]) ? {1'b1,7'd105} :
		  (single[106])? {1'b0,7'd106} : (double[106]) ? {1'b1,7'd106} :
		  (single[107])? {1'b0,7'd107} : (double[107]) ? {1'b1,7'd107} :
		  (single[108])? {1'b0,7'd108} : (double[108]) ? {1'b1,7'd108} :
		  (single[109])? {1'b0,7'd109} : (double[109]) ? {1'b1,7'd109} :
		  (single[110])? {1'b0,7'd110} : (double[110]) ? {1'b1,7'd110} :
		  (single[111])? {1'b0,7'd111} : (double[111]) ? {1'b1,7'd111} :
		  (single[112])? {1'b0,7'd112} : (double[112]) ? {1'b1,7'd112} :
		  (single[113])? {1'b0,7'd113} : (double[113]) ? {1'b1,7'd113} :
		  (single[114])? {1'b0,7'd114} : (double[114]) ? {1'b1,7'd114} :
		  (single[115])? {1'b0,7'd115} : (double[115]) ? {1'b1,7'd115} :
		  (single[116])? {1'b0,7'd116} : (double[116]) ? {1'b1,7'd116} :
		  (single[117])? {1'b0,7'd117} : (double[117]) ? {1'b1,7'd117} :
		  (single[118])? {1'b0,7'd118} : (double[118]) ? {1'b1,7'd118} :
		  (single[119])? {1'b0,7'd119} : (double[119]) ? {1'b1,7'd119} :
		  (single[120])? {1'b0,7'd120} : (double[120]) ? {1'b1,7'd120} :
		  (single[121])? {1'b0,7'd121} : (double[121]) ? {1'b1,7'd121} :
		  (single[122])? {1'b0,7'd122} : (double[122]) ? {1'b1,7'd122} :
		  (single[123])? {1'b0,7'd123} : (double[123]) ? {1'b1,7'd123} :
		  (single[124])? {1'b0,7'd124} : (double[124]) ? {1'b1,7'd124} :
		  (single[125])? {1'b0,7'd125} : (double[125]) ? {1'b1,7'd125} :
		  (single[126])? {1'b0,7'd126} : (double[126]) ? {1'b1,7'd126} :
		  (single[127])? {1'b0,7'd127} : (double[127]) ? {1'b1,7'd127} :
		  8'b11111111;
   
   // This gives the second hit cluster location
   assign second =	(single[127])? {1'b0,7'd127} : (double[127]) ? {1'b1,7'd126} :
		(single[126])? {1'b0,7'd126} : (double[126]) ? {1'b1,7'd125} :
		  (single[125])? {1'b0,7'd125} : (double[125]) ? {1'b1,7'd124} :
		  (single[124])? {1'b0,7'd124} : (double[124]) ? {1'b1,7'd123} :
		(single[123])? {1'b0,7'd123} : (double[123]) ? {1'b1,7'd122} :
		(single[122])? {1'b0,7'd122} : (double[122]) ? {1'b1,7'd121} :
		(single[121])? {1'b0,7'd121} : (double[121]) ? {1'b1,7'd120} :
		(single[120])? {1'b0,7'd120} : (double[120]) ? {1'b1,7'd119} :
		(single[119])? {1'b0,7'd119} : (double[119]) ? {1'b1,7'd118} :
		(single[118])? {1'b0,7'd118} : (double[118]) ? {1'b1,7'd117} :
		(single[117])? {1'b0,7'd117} : (double[117]) ? {1'b1,7'd116} :
		(single[116])? {1'b0,7'd116} : (double[116]) ? {1'b1,7'd115} :
		(single[115])? {1'b0,7'd115} : (double[115]) ? {1'b1,7'd114} :
		(single[114])? {1'b0,7'd114} : (double[114]) ? {1'b1,7'd113} :
		(single[113])? {1'b0,7'd113} : (double[113]) ? {1'b1,7'd112} :
		(single[112])? {1'b0,7'd112} : (double[112]) ? {1'b1,7'd111} :
		(single[111])? {1'b0,7'd111} : (double[111]) ? {1'b1,7'd110} :
		(single[110])? {1'b0,7'd110} : (double[110]) ? {1'b1,7'd109} :
		(single[109])? {1'b0,7'd109} : (double[109]) ? {1'b1,7'd108} :
		(single[108])? {1'b0,7'd108} : (double[108]) ? {1'b1,7'd107} :
		(single[107])? {1'b0,7'd107} : (double[107]) ? {1'b1,7'd106} :
		(single[106])? {1'b0,7'd106} : (double[106]) ? {1'b1,7'd105} :
		(single[105])? {1'b0,7'd105} : (double[105]) ? {1'b1,7'd104} :
		(single[104])? {1'b0,7'd104} : (double[104]) ? {1'b1,7'd103} :
		(single[103])? {1'b0,7'd103} : (double[103]) ? {1'b1,7'd102} :
		(single[102])? {1'b0,7'd102} : (double[102]) ? {1'b1,7'd101} :
		(single[101])? {1'b0,7'd101} : (double[101]) ? {1'b1,7'd100} :
		(single[100])? {1'b0,7'd100} : (double[100]) ? {1'b1,7'd99} :
		(single[99])? {1'b0,7'd99} : (double[99]) ? {1'b1,7'd98} :
		(single[98])? {1'b0,7'd98} : (double[98]) ? {1'b1,7'd97} :
		(single[97])? {1'b0,7'd97} : (double[97]) ? {1'b1,7'd96} :
		(single[96])? {1'b0,7'd96} : (double[96]) ? {1'b1,7'd95} :
		(single[95])? {1'b0,7'd95} : (double[95]) ? {1'b1,7'd94} :
		(single[94])? {1'b0,7'd94} : (double[94]) ? {1'b1,7'd93} :
		(single[93])? {1'b0,7'd93} : (double[93]) ? {1'b1,7'd92} :
		(single[92])? {1'b0,7'd92} : (double[92]) ? {1'b1,7'd91} :
		(single[91])? {1'b0,7'd91} : (double[91]) ? {1'b1,7'd90} :
		(single[90])? {1'b0,7'd90} : (double[90]) ? {1'b1,7'd89} :
		(single[89])? {1'b0,7'd89} : (double[89]) ? {1'b1,7'd88} :
		(single[88])? {1'b0,7'd88} : (double[88]) ? {1'b1,7'd87} :
		(single[87])? {1'b0,7'd87} : (double[87]) ? {1'b1,7'd86} :
		(single[86])? {1'b0,7'd86} : (double[86]) ? {1'b1,7'd85} :
		(single[85])? {1'b0,7'd85} : (double[85]) ? {1'b1,7'd84} :
		(single[84])? {1'b0,7'd84} : (double[84]) ? {1'b1,7'd83} :
		(single[83])? {1'b0,7'd83} : (double[83]) ? {1'b1,7'd82} :
		(single[82])? {1'b0,7'd82} : (double[82]) ? {1'b1,7'd81} :
		(single[81])? {1'b0,7'd81} : (double[81]) ? {1'b1,7'd80} :
		(single[80])? {1'b0,7'd80} : (double[80]) ? {1'b1,7'd79} :
		(single[79])? {1'b0,7'd79} : (double[79]) ? {1'b1,7'd78} :
		(single[78])? {1'b0,7'd78} : (double[78]) ? {1'b1,7'd77} :
		(single[77])? {1'b0,7'd77} : (double[77]) ? {1'b1,7'd76} :
		(single[76])? {1'b0,7'd76} : (double[76]) ? {1'b1,7'd75} :
		(single[75])? {1'b0,7'd75} : (double[75]) ? {1'b1,7'd74} :
		(single[74])? {1'b0,7'd74} : (double[74]) ? {1'b1,7'd73} :
		(single[73])? {1'b0,7'd73} : (double[73]) ? {1'b1,7'd72} :
		(single[72])? {1'b0,7'd72} : (double[72]) ? {1'b1,7'd71} :
		(single[71])? {1'b0,7'd71} : (double[71]) ? {1'b1,7'd70} :
		(single[70])? {1'b0,7'd70} : (double[70]) ? {1'b1,7'd69} :
		(single[69])? {1'b0,7'd69} : (double[69]) ? {1'b1,7'd68} :
		(single[68])? {1'b0,7'd68} : (double[68]) ? {1'b1,7'd67} :
		(single[67])? {1'b0,7'd67} : (double[67]) ? {1'b1,7'd66} :
		(single[66])? {1'b0,7'd66} : (double[66]) ? {1'b1,7'd65} :
		(single[65])? {1'b0,7'd65} : (double[65]) ? {1'b1,7'd64} :
		(single[64])? {1'b0,7'd64} : (double[64]) ? {1'b1,7'd63} :
		(single[63])? {1'b0,7'd63} : (double[63]) ? {1'b1,7'd62} :
		(single[62])? {1'b0,7'd62} : (double[62]) ? {1'b1,7'd61} :
		(single[61])? {1'b0,7'd61} : (double[61]) ? {1'b1,7'd60} :
		(single[60])? {1'b0,7'd60} : (double[60]) ? {1'b1,7'd59} :
		(single[59])? {1'b0,7'd59} : (double[59]) ? {1'b1,7'd58} :
		(single[58])? {1'b0,7'd58} : (double[58]) ? {1'b1,7'd57} :
		(single[57])? {1'b0,7'd57} : (double[57]) ? {1'b1,7'd56} :
		(single[56])? {1'b0,7'd56} : (double[56]) ? {1'b1,7'd55} :
		(single[55])? {1'b0,7'd55} : (double[55]) ? {1'b1,7'd54} :
		(single[54])? {1'b0,7'd54} : (double[54]) ? {1'b1,7'd53} :
		(single[53])? {1'b0,7'd53} : (double[53]) ? {1'b1,7'd52} :
		(single[52])? {1'b0,7'd52} : (double[52]) ? {1'b1,7'd51} :
		(single[51])? {1'b0,7'd51} : (double[51]) ? {1'b1,7'd50} :
		(single[50])? {1'b0,7'd50} : (double[50]) ? {1'b1,7'd49} :
		(single[49])? {1'b0,7'd49} : (double[49]) ? {1'b1,7'd48} :
		(single[48])? {1'b0,7'd48} : (double[48]) ? {1'b1,7'd47} :
		(single[47])? {1'b0,7'd47} : (double[47]) ? {1'b1,7'd46} :
		(single[46])? {1'b0,7'd46} : (double[46]) ? {1'b1,7'd45} :
		(single[45])? {1'b0,7'd45} : (double[45]) ? {1'b1,7'd44} :
		(single[44])? {1'b0,7'd44} : (double[44]) ? {1'b1,7'd43} :
		(single[43])? {1'b0,7'd43} : (double[43]) ? {1'b1,7'd42} :
		(single[42])? {1'b0,7'd42} : (double[42]) ? {1'b1,7'd41} :
		(single[41])? {1'b0,7'd41} : (double[41]) ? {1'b1,7'd40} :
		(single[40])? {1'b0,7'd40} : (double[40]) ? {1'b1,7'd39} :
		(single[39])? {1'b0,7'd39} : (double[39]) ? {1'b1,7'd38} :
		(single[38])? {1'b0,7'd38} : (double[38]) ? {1'b1,7'd37} :
		(single[37])? {1'b0,7'd37} : (double[37]) ? {1'b1,7'd36} :
		(single[36])? {1'b0,7'd36} : (double[36]) ? {1'b1,7'd35} :
		(single[35])? {1'b0,7'd35} : (double[35]) ? {1'b1,7'd34} :
		(single[34])? {1'b0,7'd34} : (double[34]) ? {1'b1,7'd33} :
		(single[33])? {1'b0,7'd33} : (double[33]) ? {1'b1,7'd32} :
		(single[32])? {1'b0,7'd32} : (double[32]) ? {1'b1,7'd31} :
		(single[31])? {1'b0,7'd31} : (double[31]) ? {1'b1,7'd30} :
		(single[30])? {1'b0,7'd30} : (double[30]) ? {1'b1,7'd29} :
		(single[29])? {1'b0,7'd29} : (double[29]) ? {1'b1,7'd28} :
		(single[28])? {1'b0,7'd28} : (double[28]) ? {1'b1,7'd27} :
		(single[27])? {1'b0,7'd27} : (double[27]) ? {1'b1,7'd26} :
		(single[26])? {1'b0,7'd26} : (double[26]) ? {1'b1,7'd25} :
		(single[25])? {1'b0,7'd25} : (double[25]) ? {1'b1,7'd24} :
		(single[24])? {1'b0,7'd24} : (double[24]) ? {1'b1,7'd23} :
		(single[23])? {1'b0,7'd23} : (double[23]) ? {1'b1,7'd22} :
		(single[22])? {1'b0,7'd22} : (double[22]) ? {1'b1,7'd21} :
		(single[21])? {1'b0,7'd21} : (double[21]) ? {1'b1,7'd20} :
		(single[20])? {1'b0,7'd20} : (double[20]) ? {1'b1,7'd19} :
		(single[19])? {1'b0,7'd19} : (double[19]) ? {1'b1,7'd18} :
		(single[18])? {1'b0,7'd18} : (double[18]) ? {1'b1,7'd17} :
		(single[17])? {1'b0,7'd17} : (double[17]) ? {1'b1,7'd16} :
		(single[16])? {1'b0,7'd16} : (double[16]) ? {1'b1,7'd15} :
		(single[15])? {1'b0,7'd15} : (double[15]) ? {1'b1,7'd14} :
		(single[14])? {1'b0,7'd14} : (double[14]) ? {1'b1,7'd13} :
		(single[13])? {1'b0,7'd13} : (double[13]) ? {1'b1,7'd12} :
		(single[12])? {1'b0,7'd12} : (double[12]) ? {1'b1,7'd11} :
		(single[11])? {1'b0,7'd11} : (double[11]) ? {1'b1,7'd10} :
		(single[10])? {1'b0,7'd10} : (double[10]) ? {1'b1,7'd9} :
		(single[9])? {1'b0,7'd9} : (double[9]) ? {1'b1,7'd8} :
		(single[8])? {1'b0,7'd8} : (double[8]) ? {1'b1,7'd7} :
		(single[7])? {1'b0,7'd7} : (double[7]) ? {1'b1,7'd6} :
		(single[6])? {1'b0,7'd6} : (double[6]) ? {1'b1,7'd5} :
		(single[5])? {1'b0,7'd5} : (double[5]) ? {1'b1,7'd4} :
		(single[4])? {1'b0,7'd4} : (double[4]) ? {1'b1,7'd3} :
		(single[3])? {1'b0,7'd3} : (double[3]) ? {1'b1,7'd2} :
		(single[2])? {1'b0,7'd2} : (double[2]) ? {1'b1,7'd1} :
		(single[1])? {1'b0,7'd1} : (double[1]) ? {1'b1,7'd0} :
		(single[0])? {1'b0,7'd0} : 8'b11111111;
						
assign firsttemp = first[6:0];

// generate the mask based on the first hit location

assign mask = 	(firsttemp == 7'd0)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100: (firsttemp == 7'd1) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001:
		(firsttemp == 7'd2)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011: (firsttemp == 7'd3) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111:
		(firsttemp == 7'd4)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111: (firsttemp == 7'd5) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111:
		(firsttemp == 7'd6)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111: (firsttemp == 7'd7) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111:
		(firsttemp == 7'd8)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111: (firsttemp == 7'd9) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111:
		(firsttemp == 7'd10)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111: (firsttemp == 7'd11) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111:
		(firsttemp == 7'd12)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111: (firsttemp == 7'd13) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111:
		(firsttemp == 7'd14)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111: (firsttemp == 7'd15) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111:
		(firsttemp == 7'd16)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111: (firsttemp == 7'd17) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111:
		(firsttemp == 7'd18)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111: (firsttemp == 7'd19) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111:
		(firsttemp == 7'd20)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111: (firsttemp == 7'd21) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111:
		(firsttemp == 7'd22)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111: (firsttemp == 7'd23) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111:
		(firsttemp == 7'd24)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111: (firsttemp == 7'd25) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111:
		(firsttemp == 7'd26)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111: (firsttemp == 7'd27) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111:
		(firsttemp == 7'd28)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111: (firsttemp == 7'd29) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111:
		(firsttemp == 7'd30)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111: (firsttemp == 7'd31) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111:
		(firsttemp == 7'd32)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111: (firsttemp == 7'd33) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111:
		(firsttemp == 7'd34)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111: (firsttemp == 7'd35) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111:
		(firsttemp == 7'd36)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111: (firsttemp == 7'd37) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111:
		(firsttemp == 7'd38)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111: (firsttemp == 7'd39) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111:
		(firsttemp == 7'd40)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111: (firsttemp == 7'd41) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111:
		(firsttemp == 7'd42)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111: (firsttemp == 7'd43) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111:
		(firsttemp == 7'd44)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111: (firsttemp == 7'd45) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111:
		(firsttemp == 7'd46)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111: (firsttemp == 7'd47) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111:
		(firsttemp == 7'd48)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111: (firsttemp == 7'd49) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd50)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111: (firsttemp == 7'd51) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd52)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111: (firsttemp == 7'd53) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd54)? 128'b11111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd55) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd56)? 128'b11111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd57) ? 128'b11111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd58)? 128'b11111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd59) ? 128'b11111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd60)? 128'b11111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd61) ? 128'b11111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd62)? 128'b11111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd63) ? 128'b11111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd64)? 128'b11111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd65) ? 128'b11111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd66)? 128'b11111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd67) ? 128'b11111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd68)? 128'b11111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd69) ? 128'b11111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd70)? 128'b11111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd71) ? 128'b11111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd72)? 128'b11111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd73) ? 128'b11111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd74)? 128'b11111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd75) ? 128'b11111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd76)? 128'b11111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd77) ? 128'b11111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd78)? 128'b11111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd79) ? 128'b11111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd80)? 128'b11111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd81) ? 128'b11111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd82)? 128'b11111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd83) ? 128'b11111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd84)? 128'b11111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd85) ? 128'b11111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd86)? 128'b11111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd87) ? 128'b11111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd88)? 128'b11111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd89) ? 128'b11111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd90)? 128'b11111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd91) ? 128'b11111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd92)? 128'b11111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd93) ? 128'b11111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd94)? 128'b11111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd95) ? 128'b11111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd96)? 128'b11111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd97) ? 128'b11111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd98)? 128'b11111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd99) ? 128'b11111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd100)? 128'b11111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd101) ? 128'b11111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd102)? 128'b11111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd103) ? 128'b11111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd104)? 128'b11111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd105) ? 128'b11111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd106)? 128'b11111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd107) ? 128'b11111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd108)? 128'b11111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd109) ? 128'b11111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd110)? 128'b11111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd111) ? 128'b11111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd112)? 128'b11111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd113) ? 128'b11111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd114)? 128'b11111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd115) ? 128'b11111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd116)? 128'b11111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd117) ? 128'b11111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd118)? 128'b11111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd119) ? 128'b11111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd120)? 128'b11111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd121) ? 128'b11111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd122)? 128'b11110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd123) ? 128'b11100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd124)? 128'b11001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd125) ? 128'b10011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		(firsttemp == 7'd126)? 128'b00111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111: (firsttemp == 7'd127) ? 128'b01111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111:
		128'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

// the datatemp masks the first hit
//assign datatemp = data & mask;

// third hit in the data where 1st hit is masked
assign third = (datatemp[0])?7'd0:
	       (datatemp[1])?7'd1:
	       (datatemp[2])?7'd2:
	       (datatemp[3])?7'd3:
	       (datatemp[4])?7'd4:
	       (datatemp[5])?7'd5:
	       (datatemp[6])?7'd6:
	       (datatemp[7])?7'd7:
	       (datatemp[8])?7'd8:
	       (datatemp[9])?7'd9:
	       (datatemp[10])?7'd10:
	       (datatemp[11])?7'd11:
	       (datatemp[12])?7'd12:
	       (datatemp[13])?7'd13:
	       (datatemp[14])?7'd14:
	       (datatemp[15])?7'd15:
	       (datatemp[16])?7'd16:
	       (datatemp[17])?7'd17:
	       (datatemp[18])?7'd18:
	       (datatemp[19])?7'd19:
	       (datatemp[20])?7'd20:
	       (datatemp[21])?7'd21:
	       (datatemp[22])?7'd22:
	       (datatemp[23])?7'd23:
	       (datatemp[24])?7'd24:
	       (datatemp[25])?7'd25:
	       (datatemp[26])?7'd26:
	       (datatemp[27])?7'd27:
	       (datatemp[28])?7'd28:
	       (datatemp[29])?7'd29:
	       (datatemp[30])?7'd30:
	       (datatemp[31])?7'd31:
	       (datatemp[32])?7'd32:
	       (datatemp[33])?7'd33:
	       (datatemp[34])?7'd34:
	       (datatemp[35])?7'd35:
	       (datatemp[36])?7'd36:
	       (datatemp[37])?7'd37:
	       (datatemp[38])?7'd38:
	       (datatemp[39])?7'd39:
	       (datatemp[40])?7'd40:
	       (datatemp[41])?7'd41:
	       (datatemp[42])?7'd42:
	       (datatemp[43])?7'd43:
	       (datatemp[44])?7'd44:
	       (datatemp[45])?7'd45:
	       (datatemp[46])?7'd46:
	       (datatemp[47])?7'd47:
	       (datatemp[48])?7'd48:
	       (datatemp[49])?7'd49:
	       (datatemp[50])?7'd50:
	       (datatemp[51])?7'd51:
	       (datatemp[52])?7'd52:
	       (datatemp[53])?7'd53:
	       (datatemp[54])?7'd54:
	       (datatemp[55])?7'd55:
	       (datatemp[56])?7'd56:
	       (datatemp[57])?7'd57:
	       (datatemp[58])?7'd58:
	       (datatemp[59])?7'd59:
	       (datatemp[60])?7'd60:
	       (datatemp[61])?7'd61:
	       (datatemp[62])?7'd62:
	       (datatemp[63])?7'd63:
	       (datatemp[64])?7'd64:
	       (datatemp[65])?7'd65:
	       (datatemp[66])?7'd66:
	       (datatemp[67])?7'd67:
	       (datatemp[68])?7'd68:
	       (datatemp[69])?7'd69:
	       (datatemp[70])?7'd70:
	       (datatemp[71])?7'd71:
	       (datatemp[72])?7'd72:
	       (datatemp[73])?7'd73:
	       (datatemp[74])?7'd74:
	       (datatemp[75])?7'd75:
	       (datatemp[76])?7'd76:
	       (datatemp[77])?7'd77:
	       (datatemp[78])?7'd78:
	       (datatemp[79])?7'd79:
	       (datatemp[80])?7'd80:
	       (datatemp[81])?7'd81:
	       (datatemp[82])?7'd82:
	       (datatemp[83])?7'd83:
	       (datatemp[84])?7'd84:
	       (datatemp[85])?7'd85:
	       (datatemp[86])?7'd86:
	       (datatemp[87])?7'd87:
	       (datatemp[88])?7'd88:
	       (datatemp[89])?7'd89:
	       (datatemp[90])?7'd90:
	       (datatemp[91])?7'd91:
	       (datatemp[92])?7'd92:
	       (datatemp[93])?7'd93:
	       (datatemp[94])?7'd94:
	       (datatemp[95])?7'd95:
	       (datatemp[96])?7'd96:
	       (datatemp[97])?7'd97:
	       (datatemp[98])?7'd98:
               (datatemp[99])?7'd99:
	       (datatemp[100])?7'd100:
	       (datatemp[101])?7'd101:
	       (datatemp[102])?7'd102:
	       (datatemp[103])?7'd103:
	       (datatemp[104])?7'd104:
	       (datatemp[105])?7'd105:
	       (datatemp[106])?7'd106:
               (datatemp[107])?7'd107:
	       (datatemp[108])?7'd108:
	       (datatemp[109])?7'd109:
	       (datatemp[110])?7'd110:
	       (datatemp[111])?7'd111:
	       (datatemp[112])?7'd112:
	       (datatemp[113])?7'd113:
	       (datatemp[114])?7'd114:
	       (datatemp[115])?7'd115:
	       (datatemp[116])?7'd116:
	       (datatemp[117])?7'd117:
	       (datatemp[118])?7'd118:
	       (datatemp[119])?7'd119:
	       (datatemp[120])?7'd120:
	       (datatemp[121])?7'd121:
	       (datatemp[122])?7'd122:
	       (datatemp[123])?7'd123:
	       (datatemp[124])?7'd124:
	       (datatemp[125])?7'd125:
	       (datatemp[126])?7'd126:
	       (datatemp[127])?7'd127:7'b1111111;
	       
// If the third location is same as second ,OR if there is only one hit, then enter the right address, if not enter all ones.
assign totaladdr[7:0] = (first != 8'b11111111)? first:8'b11111111;
assign totaladdr[15:8] = (second != 8'b11111111)? second:8'b11111111;

//delay delayClk (.In(BCclk),.Out(lclClk));
/* 						
always @ (negedge BCclk)
begin
	if ((third[6:0]==second[6:0])|(third[6:0]==first[6:0])|(first==second))
	  count<= 1'b0;
	else
	  count<=  1'b1;
end
 */  
endmodule
