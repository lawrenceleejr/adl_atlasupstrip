
`timescale 1ns/10ps
module cluster_mux(
	input [127:0] data_i,
	input [6:0] sel,
	output [3:0] data_o);

assign data_o = (sel==127)?data_i[127:124]:
		(sel==126)?data_i[126:123]:
		(sel==125)?data_i[125:122]:
		(sel==124)?data_i[124:121]:
		(sel==123)?data_i[123:120]:
		(sel==122)?data_i[122:119]:
		(sel==121)?data_i[121:118]:
		(sel==120)?data_i[120:117]:
		(sel==119)?data_i[119:116]:
		(sel==118)?data_i[118:115]:
		(sel==117)?data_i[117:114]:
		(sel==116)?data_i[116:113]:
		(sel==115)?data_i[115:112]:
		(sel==114)?data_i[114:111]:
		(sel==113)?data_i[113:110]:
		(sel==112)?data_i[112:109]:
		(sel==111)?data_i[111:108]:
		(sel==110)?data_i[110:107]:
		(sel==109)?data_i[109:106]:
		(sel==108)?data_i[108:105]:
		(sel==107)?data_i[107:104]:
		(sel==106)?data_i[106:103]:
		(sel==105)?data_i[105:102]:
		(sel==104)?data_i[104:101]:
		(sel==103)?data_i[103:100]:
		(sel==102)?data_i[102:99]:
		(sel==101)?data_i[101:98]:
		(sel==100)?data_i[100:97]:
		(sel==99)?data_i[99:96]:
		(sel==98)?data_i[98:95]:
		(sel==97)?data_i[97:94]:
		(sel==96)?data_i[96:93]:
		(sel==95)?data_i[95:92]:
		(sel==94)?data_i[94:91]:
		(sel==93)?data_i[93:90]:
		(sel==92)?data_i[92:89]:
		(sel==91)?data_i[91:88]:
		(sel==90)?data_i[90:87]:
		(sel==89)?data_i[89:86]:
		(sel==88)?data_i[88:85]:
		(sel==87)?data_i[87:84]:
		(sel==86)?data_i[86:83]:
		(sel==85)?data_i[85:82]:
		(sel==84)?data_i[84:81]:
		(sel==83)?data_i[83:80]:
		(sel==82)?data_i[82:79]:
		(sel==81)?data_i[81:78]:
		(sel==80)?data_i[80:77]:
		(sel==79)?data_i[79:76]:
		(sel==78)?data_i[78:75]:
		(sel==77)?data_i[77:74]:
		(sel==76)?data_i[76:73]:
		(sel==75)?data_i[75:72]:
		(sel==74)?data_i[74:71]:
		(sel==73)?data_i[73:70]:
		(sel==72)?data_i[72:69]:
		(sel==71)?data_i[71:68]:
		(sel==70)?data_i[70:67]:
		(sel==69)?data_i[69:66]:
		(sel==68)?data_i[68:65]:
		(sel==67)?data_i[67:64]:
		(sel==66)?data_i[66:63]:
		(sel==65)?data_i[65:62]:
		(sel==64)?data_i[64:61]:
		(sel==63)?data_i[63:60]:
		(sel==62)?data_i[62:59]:
		(sel==61)?data_i[61:58]:
		(sel==60)?data_i[60:57]:
		(sel==59)?data_i[59:56]:
		(sel==58)?data_i[58:55]:
		(sel==57)?data_i[57:54]:
		(sel==56)?data_i[56:53]:
		(sel==55)?data_i[55:52]:
		(sel==54)?data_i[54:51]:
		(sel==53)?data_i[53:50]:
		(sel==52)?data_i[52:49]:
		(sel==51)?data_i[51:48]:
		(sel==50)?data_i[50:47]:
		(sel==49)?data_i[49:46]:
		(sel==48)?data_i[48:45]:
		(sel==47)?data_i[47:44]:
		(sel==46)?data_i[46:43]:
		(sel==45)?data_i[45:42]:
		(sel==44)?data_i[44:41]:
		(sel==43)?data_i[43:40]:
		(sel==42)?data_i[42:39]:
		(sel==41)?data_i[41:38]:
		(sel==40)?data_i[40:37]:
		(sel==39)?data_i[39:36]:
		(sel==38)?data_i[38:35]:
		(sel==37)?data_i[37:34]:
		(sel==36)?data_i[36:33]:
		(sel==35)?data_i[35:32]:
		(sel==34)?data_i[34:31]:
		(sel==33)?data_i[33:30]:
		(sel==32)?data_i[32:29]:
		(sel==31)?data_i[31:28]:
		(sel==30)?data_i[30:27]:
		(sel==29)?data_i[29:26]:
		(sel==28)?data_i[28:25]:
		(sel==27)?data_i[27:24]:
		(sel==26)?data_i[26:23]:
		(sel==25)?data_i[25:22]:
		(sel==24)?data_i[24:21]:
		(sel==23)?data_i[23:20]:
		(sel==22)?data_i[22:19]:
		(sel==21)?data_i[21:18]:
		(sel==20)?data_i[20:17]:
		(sel==19)?data_i[19:16]:
		(sel==18)?data_i[18:15]:
		(sel==17)?data_i[17:14]:
		(sel==16)?data_i[16:13]:
		(sel==15)?data_i[15:12]:
		(sel==14)?data_i[14:11]:
		(sel==13)?data_i[13:10]:
		(sel==12)?data_i[12:9]:
		(sel==11)?data_i[11:8]:
		(sel==10)?data_i[10:7]:
		(sel==9)?data_i[9:6]:
		(sel==8)?data_i[8:5]:
		(sel==7)?data_i[7:4]:
		(sel==6)?data_i[6:3]:
		(sel==5)?data_i[5:2]:
		(sel==4)?data_i[4:1]:
		(sel==3)?data_i[3:0]:
		(sel==2)?{data_i[2:0],1'b0}:
		(sel==1)?{data_i[1:0],2'b0}:
		(sel==0)?{data_i[0],3'b0}:4'b0;
endmodule
