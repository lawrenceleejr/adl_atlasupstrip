-------------------------------------------------------------------------------
-- Title         : OSRAM SCDV5540 Display Controller Characters
-- Project       : General Purpose Core
-------------------------------------------------------------------------------
-- File          : DisplayCharacters.vhd
-- Author        : Ryan Herbst, rherbst@slac.stanford.edu
-- Created       : 12/06/2007
-------------------------------------------------------------------------------
-- Description:
-- Package for display chracter lookup table.
-------------------------------------------------------------------------------
-- Copyright (c) 2007 by Ryan Herbst. All rights reserved.
-------------------------------------------------------------------------------
-- Modification history:
-- 12/06/2007: created.
-------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

package DisplayCharacters is

   -- Types For Character Lookup
   subtype DISPCHAR  is STD_LOGIC_VECTOR(24 downto 0);
   type    DISPTABLE is array ( NATURAL range <> ) of DISPCHAR;

   -- Constants For Charactors
   constant DISPMAX    : natural   := 18;
   constant DISPLOOKUP : DISPTABLE := (
         0 => "01110" & -- Hex 0
              "10011" &
              "10101" &
              "11001" &
              "01110",
         1 => "00100" & -- Hex 1
              "01100" &
              "00100" &
              "00100" &
              "11111",
         2 => "11110" & -- Hex 2
              "00001" &
              "00110" &
              "01000" &
              "11111",
         3 => "11110" & -- Hex 3
              "00001" &
              "01110" &
              "00001" &
              "11110",
         4 => "00110" & -- Hex 4
              "01010" &
              "11111" &
              "00010" &
              "00010",
         5 => "11111" & -- Hex 5
              "10000" &
              "11110" &
              "00001" &
              "11110",
         6 => "00110" & -- Hex 6
              "01000" &
              "11110" &
              "10001" &
              "01110",
         7 => "11111" & -- Hex 7
              "00010" &
              "00100" &
              "01000" &
              "01000",
         8 => "01110" & -- Hex 8
              "10001" &
              "01110" &
              "10001" &
              "01110",
         9 => "01110" & -- Hex 9
              "10001" &
              "01111" &
              "00010" &
              "01100",
        10 => "00100" & -- Hex A
              "01010" &
              "11111" &
              "10001" &
              "10001",
        11 => "11110" & -- Hex B
              "01001" &
              "01110" &
              "01001" &
              "11110",
        12 => "01111" & -- Hex C
              "10000" &
              "10000" &
              "10000" &
              "11111",
        13 => "11110" & -- Hex D
              "01001" &
              "01001" &
              "01001" &
              "11110",
        14 => "11111" & -- Hex E
              "10000" &
              "11111" &
              "10000" &
              "11111",
        15 => "11111" & -- Hex F
              "10000" &
              "11110" &
              "10000" &
              "10000",
        16 => "11110" & -- State P = No PLL Lock
              "10001" &
              "11110" &
              "10000" &
              "10000",
        17 => "10001" & -- State N = No Link
              "11001" &
              "10101" &
              "10011" &
              "10001",
        18 => "10000" & -- State L = Link
              "10000" &
              "10000" &
              "10000" &
              "11111" 
   );

end DisplayCharacters;
